`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:38:25 02/27/2013 
// Design Name: 
// Module Name:    operation 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module operation(
	input clk_100MHz,
	input operation_enable,
	input [7:0] data_in,
	output [7:0] data_out);
endmodule
